`timescale 1ns / 1ps
//Subject:     CO project 4 - Pipe CPU 1
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------
module Pipe_CPU_1(
    clk_i,
    rst_i
);
    
/****************************************
I/O ports
****************************************/
input clk_i;
input rst_i;

/****************************************
Internal signal
****************************************/
/**** IF stage ****/
wire [31:0]	pc_next_IF, pc_in_IF, pc_out_IF, instr_IF;

/**** ID stage ****/
wire [31:0]	pc_next_ID, instr_ID, RSdata_ID, RTdata_ID, extended_ID;

//control signal
wire 		RegWrite_ID, ALUSrc_ID, RegDst_ID, Branch_ID, MemRead_ID, MemWrite_ID, MemtoReg_ID;
wire [1:0]  BranchType_ID;
wire [2:0]	ALU_op_ID;

/**** EX stage ****/
wire [31:0]	pc_next_EX, RSdata_EX, RTdata_EX, extended_EX, shifted_EX, selected_EX, result_EX, pc_branch_EX, ALUSource1_EX, MuxB_o, ALUSource2_EX;
wire [4:0]	Src_EX, Dst0_EX, Dst1_EX, RDaddr_EX;

//control signal
wire [4:0]  MEM_EX;
wire [3:0]	ALUCtrl_EX;
wire [2:0]	ALU_op_EX;
wire [1:0]	WB_EX;
wire [1:0]  BranchType_EX;
wire		    RegDst_EX, ALUSrc_EX, zero_EX;
wire        Forward_A, Forward_B;

/**** MEM stage ****/
wire [31:0]	pc_branch_MEM, result_MEM, RTdata_MEM, Memdata_MEM;
wire [4:0]	RDaddr_MEM;

//control signal
wire [1:0]	WB_MEM;
wire 		Branch_MEM, MemRead_MEM, MemWrite_MEM, zero_MEM;
wire        PCSrc_MEM, Bch_MEM;

/**** WB stage ****/
wire [31:0]	RDdata_WB, Memdata_WB, result_WB;
wire [4:0]	RDaddr_WB;

//control signal
wire 		RegWrite_WB, MemtoReg_WB;

wire        PC_Write;
wire			IF_ID_Write;
wire        IF_Flush;
wire        ID_Flush;
wire        EX_Flush;
/****************************************
Instantiate modules
****************************************/
//Instantiate the components in IF stage
MUX_2to1 #(.size(32)) Mux0(
	.data0_i(pc_next_IF),
	.data1_i(pc_branch_MEM),
	.select_i(PCSrc_MEM),
	.data_o(pc_in_IF)
);

ProgramCounter PC(
	.clk_i(clk_i),
	.rst_i(rst_i),
	.pc_write(PC_Write),
	.pc_in_i(pc_in_IF),
	.pc_out_o(pc_out_IF)
);

Instruction_Memory IM(
	.addr_i(pc_out_IF),
	.instr_o(instr_IF)
);
			
Adder Add_pc(
	.src1_i(pc_out_IF),
	.src2_i(32'd4),
	.sum_o(pc_next_IF)
);

Pipe_Reg #(.size(64)) IF_ID(
	.clk_i(clk_i),
	.rst_i(rst_i),
	.write(IF_ID_Write),
	.flush(IF_Flush),
	.data_i({pc_next_IF, instr_IF}),
	.data_o({pc_next_ID, instr_ID})
);

//Instantiate the components in ID stage
Reg_File RF(
	.clk_i(clk_i),
	.rst_i(rst_i),
	.RSaddr_i(instr_ID[25:21]),
	.RTaddr_i(instr_ID[20:16]),
	.RDaddr_i(RDaddr_WB),
	.RDdata_i(RDdata_WB),
	.RegWrite_i(RegWrite_WB),
	.RSdata_o(RSdata_ID),
	.RTdata_o(RTdata_ID)
);

Decoder Control(
	.instr_op_i(instr_ID[31:26]),
	.RegWrite_o(RegWrite_ID),
	.ALU_op_o(ALU_op_ID),
	.ALUSrc_o(ALUSrc_ID),
	.RegDst_o(RegDst_ID),
	.Branch_o(Branch_ID),
	.BranchType_o(BranchType_ID),
	.MemRead_o(MemRead_ID),
	.MemWrite_o(MemWrite_ID),
	.MemtoReg_o(MemtoReg_ID)
);

HazardDetection HazardDetection(
	.EX_MemRead(MEM_EX[3]), // MemRead_EX
	.EX_Rt(Dst0_EX),
	.ID_Rs(instr_ID[25:21]),
	.ID_Rt(instr_ID[20:16]),
	.PCSrc(PCSrc_MEM),
	.PC_Write(PC_Write),
	.IF_ID_Write(IF_ID_Write),
	.IF_Flush(IF_Flush),
	.ID_Flush(ID_Flush),
	.EX_Flush(EX_Flush)
);

Sign_Extend Sign_Extend(
	.data_i(instr_ID[15:0]),
	.data_o(extended_ID)
);	

Pipe_Reg #(.size(64)) ID_EX_ReadData(
	.clk_i(clk_i),
    .rst_i(rst_i),
	.write(1'b1),
	.flush(1'b0),
    .data_i({RSdata_ID,RTdata_ID}),
    .data_o({RSdata_EX,RTdata_EX})
);

Pipe_Reg #(.size(12)) ID_EX_Control(
	.clk_i(clk_i),
    .rst_i(rst_i),
	.write(1'b1),
	.flush(ID_Flush),
    .data_i({RegWrite_ID, MemtoReg_ID, Branch_ID, BranchType_ID, MemRead_ID, MemWrite_ID, RegDst_ID, ALU_op_ID, ALUSrc_ID}),
    .data_o({WB_EX, MEM_EX, RegDst_EX, ALU_op_EX, ALUSrc_EX})
);

Pipe_Reg #(.size(32)) ID_EX_PC_Add4(
	.clk_i(clk_i),
    .rst_i(rst_i),
	.write(1'b1),
	.flush(1'b0),
    .data_i(pc_next_ID),
    .data_o(pc_next_EX)
);

Pipe_Reg #(.size(32)) ID_EX_Instruction_Extended(
	.clk_i(clk_i),
    .rst_i(rst_i),
	.write(1'b1),
	.flush(1'b0),
    .data_i(extended_ID),
    .data_o(extended_EX)
);


Pipe_Reg #(.size(15)) ID_EX_Instruction(
	.clk_i(clk_i),
    .rst_i(rst_i),
	.write(1'b1),
	.flush(1'b0),
    .data_i(instr_ID[25:11]),
    .data_o({Src_EX, Dst0_EX, Dst1_EX})
);

//Instantiate the components in EX stage	   
Shift_Left_Two_32 Shifter(
	.data_i(extended_EX),
	.data_o(shifted_EX)
);

Forwarding Forwarding_Unit(
	.EX_Rs(Src_EX),
	.EX_Rt(Dst0_EX),
	.MEM_Rd(RDadddr_MEM),
	.MEM_RegWrite(WB_MEM[0]), //RegWrite_MEM
	.WB_Rd(RDaddr_WB),
	.WB_RegWrite(RegWrite_WB),
	.Forward_A(Forward_A),
	.Forward_B(Forward_B)
    );

MUX_3to1 #(.size(32)) MuxA(
	.data0_i(RSdata_EX),
	.data1_i(result_MEM),
	.data2_i(RDdata_WB),
	.select_i(Forward_A),
    .data_o(ALUSource1_EX)
);

MUX_3to1 #(.size(32)) MuxB(
	.data0_i(RTdata_EX),
	.data1_i(result_MEM),
	.data2_i(RDdata_WB),
	.select_i(Forward_B),
    .data_o(MuxB_o)
);


MUX_2to1 #(.size(32)) Mux_ALU_Source2(
	.data0_i(MuxB_o),
	.data1_i(extended_EX),
	.select_i(ALUSrc_EX),
    .data_o(ALUSource2_EX)
);

ALU ALU(
	.src1_i(ALUSource1_EX),
	.src2_i(ALUSource2_EX),
	.ctrl_i(ALUCtrl_EX),
	.result_o(result_EX),
	.zero_o(zero_EX)
);
		
ALU_Ctrl ALU_Control(
	.funct_i(extended_EX[5:0]),
	.ALUOp_i(ALU_op_EX),
	.ALUCtrl_o(ALUCtrl_EX)
);

MUX_2to1 #(.size(5)) Mux2(
	.data0_i(Dst0_EX),
	.data1_i(Dst1_EX),
	.select_i(RegDst_EX),
    .data_o(RDaddr_EX)
);

Adder Add_pc_branch(
	.src1_i(pc_next_EX),
	.src2_i(shifted_EX),
	.sum_o(pc_branch_EX)
);

Pipe_Reg #(.size(7)) EX_MEM_Control(
	.clk_i(clk_i),
        .rst_i(rst_i),
	.write(1'b1),
	.flush(EX_Flush),
        .data_i({WB_EX, MEM_EX}),
        .data_o({WB_MEM, Branch_MEM, BranchType_MEM, MemRead_MEM, MemWrite_MEM})
);

Pipe_Reg #(.size(129)) EX_MEM_data(
	.clk_i(clk_i),
        .rst_i(rst_i),
	.write(1'b1),
	.flush(1'b0),
        .data_i({pc_branch_EX, zero_EX, result_EX, MuxB_o, RDaddr_EX}),
        .data_o({pc_branch_MEM, zero_MEM, result_MEM, RTdata_MEM, RDaddr_MEM})
);


MUX_4to1 #(.size(1)) BranchType_Mux(
	.data0_i(zero_MEM),
	.data1_i(~(zero_MEM | result_MEM[0])),
	.data2_i(~result_MEM),
	.data3_i(~zero_MEM),
	.select_i(BranchType_MEM),
    .data_o(Bch_MEM)
);

and Branch (PCSrc_MEM, Bch_MEM, Branch_MEM);

//Instantiate the components in MEM stage
Data_Memory DM(
	.clk_i(clk_i),
	.addr_i(result_MEM),
	.data_i(RTdata_MEM),
	.MemRead_i(MemRead_MEM),
	.MemWrite_i(MemWrite_MEM),
	.data_o(Memdata_MEM)
);

Pipe_Reg #(.size(71)) MEM_WB(
	.clk_i(clk_i),
	.rst_i(rst_i),
	.data_i({WB_MEM, Memdata_MEM, result_MEM, RDaddr_MEM}),
	.data_o({RegWrite_WB, MemtoReg_WB, Memdata_WB, result_WB, RDaddr_WB})
);


//Instantiate the components in WB stage
MUX_2to1 #(.size(32)) Mux_WB(
	.data0_i(result_WB),
	.data1_i(Memdata_WB),
	.select_i(MemtoReg_WB),
	.data_o(RDdata_WB)
);

/****************************************
signal assignment
****************************************/

endmodule
